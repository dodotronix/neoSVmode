
module param_module #(parameter int PARAM1=20,
                      parameter int PARAM2=30,
                      parameter logic PARAM3=40)(

                      input logic a,
                      output logic b);

    // body of the param_module

endmodule
