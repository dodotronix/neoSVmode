
module io_simple_module_ansi(
    input logic clk,
    input logic en,
    input logic rst,
    input logic [7:0] data,
    output logic res1,
    output logic res2,
    output logic fdbk);

    // body of the io_module

endmodule
