
module interface_module_ansi (
    t_clock.consumer Clk_x,
    t_bus.master bus_x,
    iface.general general_x,
    t_control.consumer ctrl_x, 
    input c,
    output d
    );

    // bodu of the interface_module_ansi 

endmodule
